/*

Copyright (C) 2012

Arvind <arvind@csail.mit.edu>
Muralidaran Vijayaraghavan <vmurali@csail.mit.edu>

Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

*/

import Vector::*;

typedef 32 AddrSz;
typedef Bit#(AddrSz) Addr;

typedef 32 DataSz;
typedef Bit#(DataSz) Data;

typedef Bit#(8) Byte;
typedef Bit#(16) Word;
typedef Bit#(32) LongWord;

typedef union tagged {
    Byte Byte;
    Word Word;
} Number deriving (Bits, Eq, FShow);

instance Literal#(Number);
    function Number fromInteger (Integer x);
        return tagged Word fromInteger(x);
    endfunction
    function Bool inLiteralRange(Number target, Integer i);
        if (target matches tagged Word .w &&& fromInteger(i) >= 256)
            return False;
        else if (target matches tagged Word .w &&& fromInteger(i) >= 65536)
            return False;
        else
            return True;
    endfunction
endinstance

instance Arith#(Number);
    function Number \+ (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word + y.Word);
        else
            ret = tagged Byte (x.Byte + y.Byte);
        return ret;
    endfunction
    function Number \- (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word - y.Word);
        else
            ret = tagged Byte (x.Byte - y.Byte);
        return ret;
    endfunction
    function Number negate (Number x);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (-x.Word);
        else
            ret = tagged Byte (-x.Byte);
        return ret;
    endfunction
    function Number \* (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word * y.Word);
        else
            ret = tagged Byte (x.Byte * y.Byte);
        return ret;
    endfunction
    function Number \/ (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word / y.Word);
        else
            ret = tagged Byte (x.Byte / y.Byte);
        return ret;
    endfunction
    function Number \% (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word % y.Word);
        else
            ret = tagged Byte (x.Byte % y.Byte);
        return ret;
    endfunction
endinstance

instance Bitwise#(Number);
    function Number \& (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word & y.Word);
        else
            ret = tagged Byte (x.Byte & y.Byte);
        return ret;
    endfunction
    function Number \| (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word | y.Word);
        else
            ret = tagged Byte (x.Byte | y.Byte);
        return ret;
    endfunction
    function Number \^ (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word ^ y.Word);
        else
            ret = tagged Byte (x.Byte ^ y.Byte);
        return ret;
    endfunction
    function Number \~^ (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word ~^ y.Word);
        else
            ret = tagged Byte (x.Byte ~^ y.Byte);
        return ret;
    endfunction
    function Number \^~ (Number x, Number y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word ^~ y.Word);
        else
            ret = tagged Byte (x.Byte ^~ y.Byte);
        return ret;
    endfunction
    function Number invert (Number x);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (~x.Word);
        else
            ret = tagged Byte (~x.Byte);
        return ret;
    endfunction
    function Number \<< (Number x, y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word << y);
        else
            ret = tagged Byte (x.Byte << y);
        return ret;
    endfunction
    function Number \>> (Number x, y);
        Number ret = ?;
        if (x matches tagged Word .w)
            ret = tagged Word (x.Word >> y);
        else
            ret = tagged Byte (x.Byte >> y);
        return ret;
    endfunction
    function Bit#(1) msb (Number x);
        Bit#(1) ret = ?;
        if (x matches tagged Word .w)
            ret = msb(x.Word);
        else
            ret = msb(x.Byte);
        return ret;
    endfunction
    function Bit#(1) lsb (Number x);
        Bit#(1) ret = ?;
        if (x matches tagged Word .w)
            ret = lsb(x.Word);
        else
            ret = lsb(x.Byte);
        return ret;
    endfunction
endinstance
