import Ehr::*;
import Vector::*;
import GetPut::*;

//////////////////
// SFifo interface 

interface SFifo#(numeric type n, type dt, type st);
    method Bool search(st x);
    method Bool notFull;
    method Action enq(dt x);
    method Action enq2(dt x, dt y);
    method Bool notEmpty;
    method Action deq;
    method Action deq2;
    method dt first;
    method Action clear;
endinterface
/*
//////////////////
// Pipeline SFIFO

// deq < search < enq < clear
module mkPipelineSFifo( function Bool isFound(dt x, st y), SFifo#(n, dt, st) ifc ) provisos (Bits#(dt,dtSz));
    // n is size of the FIFO
    // dt is data type
    // st is search type
    Vector#(n, Reg#(dt))    data     <- replicateM(mkRegU());
    Ehr#(2, Bit#(TLog#(n))) enqP     <- mkEhr(0);
    Ehr#(2, Bit#(TLog#(n))) deqP     <- mkEhr(0);
    Ehr#(3, Bool)           empty    <- mkEhr(True);
    Ehr#(3, Bool)           full     <- mkEhr(False);
    Bit#(TLog#(n))          max_index = fromInteger(valueOf(n)-1);

    method Bool search(st x);
        // look between deqP[1] and enqP[0]
        Bool ret = False;
        Bool enqP_lt_deqP = enqP[0] < deqP[1];
        for( Integer i = 0 ; i < valueOf(n) ; i = i+1 ) begin
            Bool lt_enqP = fromInteger(i) < enqP[0];
            Bool gte_deqP = fromInteger(i) >= deqP[1];
            Bool is_match = isFound(data[i], x);
            if( full[1] || (enqP_lt_deqP && lt_enqP) || (enqP_lt_deqP && gte_deqP) || (lt_enqP && gte_deqP) ) begin
                // index i is valid
                if( is_match ) begin
                    ret = True;
                end
            end
        end
        return ret;
    endmethod

    method Bool notFull = !full[1];

    method Action enq(dt x) if( !full[1] );
        data[enqP[0]] <= x;
        empty[1] <= False;
        enqP[0] <= (enqP[0] == max_index) ? 0 : enqP[0] + 1;
        if( enqP[1] == deqP[1] ) begin
            full[1] <= True;
        end
    endmethod

    method Bool notEmpty = !empty[0];

    method Action deq if( !empty[0] );
        // Tell later stages a dequeue was requested
        full[0] <= False;
        deqP[0] <= (deqP[0] == max_index) ? 0 : deqP[0] + 1;
        if( deqP[1] == enqP[0] ) begin
            empty[0] <= True;
        end
    endmethod

    method dt first if( !empty[0] );
        return data[deqP[0]];
    endmethod

    method Action clear;
        enqP[1] <= 0;
        deqP[1] <= 0;
        empty[2] <= True;
        full[2] <= False;
    endmethod
endmodule*/

////////////////
// Bypass SFIFO

module mkBypassSFifo( function Bool isFound(dt x, st y), SFifo#(n, dt, st) ifc ) provisos (Bits#(dt,dtSz));
    // n is size of fifo
    // t is data type of fifo
    Vector#(n, Ehr#(2,dt))  data     <- replicateM(mkEhr(?));
    Ehr#(2, Bit#(TLog#(n))) enqP     <- mkEhr(0);
    Ehr#(2, Bit#(TLog#(n))) deqP     <- mkEhr(0);
    Ehr#(3, Bool)           empty    <- mkEhr(True);
    Ehr#(3, Bool)           full     <- mkEhr(False);
    Bit#(TLog#(n))          max_index = fromInteger(valueOf(n)-1);

    method Bool search(st x);
        // look between deqP[0] and enqP[0]
        Bool ret = False;
        Bool enqP_lt_deqP = enqP[0] < deqP[0];
        for( Integer i = 0 ; i < valueOf(n) ; i = i+1 ) begin
            Bool lt_enqP = fromInteger(i) < enqP[0];
            Bool gte_deqP = fromInteger(i) >= deqP[0];
            Bool is_match = isFound(data[i][0], x);
            if( full[0] || (enqP_lt_deqP && lt_enqP) || (enqP_lt_deqP && gte_deqP) || (lt_enqP && gte_deqP) ) begin
                // index i is valid
                if( is_match ) begin
                    ret = True;
                end
            end
        end
        return ret;
    endmethod

    method Bool notFull = !full[0];

    method Action enq(dt x) if( !full[0] );
        data[enqP[0]][0] <= x;
        empty[0] <= False;
        enqP[0] <= (enqP[0] == max_index) ? 0 : enqP[0] + 1;
        if( enqP[1] == deqP[0] ) begin
            full[0] <= True;
        end
    endmethod

    // THIS is a dangerous method, does not check limits for full if 1 slot empty
    method Action enq2(dt x, dt y) if( !full[0] );
        data[enqP[0]][0] <= x;
        data[(enqP[0] == max_index) ? 0 : enqP[0] + 1][0] <= y;
        empty[0] <= False;
        enqP[0] <= (enqP[0] == max_index) ? 1 : ((enqP[0] == max_index - 1) ? 0 : enqP[0] + 2);
        if( enqP[1] == deqP[0] ) begin
            full[0] <= True;
        end

        $display("     Scoreboard: ENQ enqP[1]: ", fshow(enqP[1]), ", deqP[0]", fshow(deqP[0]), ", empty: ", empty[2], ", full: ", full[2]);
        $display("      0: %h", data[0][1], ", 1: %h", data[1][1], ", 2: %h", data[2][1], ", 3: %h", data[3][1], ", 4: %h", data[4][1], ", 5: %h", data[5][1], ", 6: %h", data[6][1], ", 7: %h", data[7][1], ", 8: %h", data[8][1], ", 9: %h", data[9][1], ", 10: %h", data[10][1], ", 11: %h", data[11][1], ", 12: %h", data[12][1], ", 13: %h", data[13][1]);
    endmethod

    method Bool notEmpty = !empty[1];

    method Action deq if( !empty[1] );
        // Tell later stages a dequeue was requested
        full[1] <= False;
        deqP[0] <= (deqP[0] == max_index) ? 0 : deqP[0] + 1;
        if( deqP[1] == enqP[1] ) begin
            empty[1] <= True;
        end
    endmethod

    // THIS is a dangerous method, does not check limits for empty
    method Action deq2 if( !empty[1] );
        // Tell later stages a dequeue was requested
        full[1] <= False;
        deqP[0] <= (deqP[0] == max_index) ? 1 : ((deqP[0] == max_index - 1) ? 0 : deqP[0] + 2);
        if( deqP[1] == enqP[1] ) begin
            empty[1] <= True;
        end

        $display("     Scoreboard: DEQ enqP[1]: ", fshow(enqP[1]), ", deqP[0]", fshow(deqP[1]), ", empty: ", empty[2], ", full: ", full[2]);
        $display("      0: %h", data[0][1], ", 1: %h", data[1][1], ", 2: %h", data[2][1], ", 3: %h", data[3][1], ", 4: %h", data[4][1], ", 5: %h", data[5][1], ", 6: %h", data[6][1], ", 7: %h", data[7][1], ", 8: %h", data[8][1], ", 9: %h", data[9][1], ", 10: %h", data[10][1], ", 11: %h", data[11][1], ", 12: %h", data[12][1], ", 13: %h", data[13][1]);

    endmethod

    method dt first if( !empty[1] );
        return data[deqP[0]][1];
    endmethod

    method Action clear;
        enqP[1] <= 0;
        deqP[1] <= 0;
        empty[2] <= True;
        full[2] <= False;
    endmethod
endmodule

